LIBRARY IEEE; -- THU VIEN CHUAN IEEE
USE IEEE.STD_LOGIC_1164.ALL; -- SU DUNG GOI THU VIEN HO TRO CAC PHEP TOAN LOGIC
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
-- FILE MO PHONG QUA TRINH TRUYEN NHAN CUA BO UART.
ENTITY TRANSFER IS 
PORT(
	CLK	 : IN  STD_LOGIC:='0';
	TX	 : OUT STD_LOGIC:='1';
	RX	 : IN  STD_LOGIC;
	RX_DATA	 : BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0));
END TRANSFER;

ARCHITECTURE TRANSFER_ARCH OF TRANSFER IS
SIGNAL RST_N	 : STD_LOGIC:='1';
SIGNAL PULSE	 : STD_LOGIC:='0';
SIGNAL TX_ENA	 : STD_LOGIC:='0';
SIGNAL TX_DATA	 : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL TX_BUSY	 : STD_LOGIC;
SIGNAL TX_DONE	 : STD_LOGIC;
SIGNAL RX_BUSY	 : STD_LOGIC;
SIGNAL RX_ERROR  : STD_LOGIC;
SIGNAL CNT_DATA  : STD_LOGIC_VECTOR(15 DOWNTO 0):=(OTHERS=>'0');
--
TYPE ASCII_ARRAY IS ARRAY (0 TO 5) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL HELLO : ASCII_ARRAY := (
    0 => X"48",  -- 'H'
    1 => X"45",  -- 'E'
    2 => X"4C",  -- 'L'
    3 => X"4C",  -- 'L'
    4 => X"4F",  -- 'O'
    5 => X"0A"   -- '\n' 
);
--
COMPONENT UART
    PORT (
        CLK      : IN  STD_LOGIC;
        RST_N    : IN  STD_LOGIC;
        TX_ENA   : IN  STD_LOGIC;
        TX_DATA  : IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
        TX       : OUT STD_LOGIC;
        TX_BUSY  : OUT STD_LOGIC;
        TX_DONE  : OUT STD_LOGIC;
        RX       : IN  STD_LOGIC;
        RX_BUSY  : OUT STD_LOGIC;
        RX_ERROR : OUT STD_LOGIC;
        RX_DATA  : BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END COMPONENT;
--
BEGIN
UA: UART
    PORT MAP (
        CLK      => CLK,
        RST_N    => RST_N,
        TX_ENA   => TX_ENA,
        TX_DATA  => TX_DATA,
        TX       => TX,
        TX_BUSY  => TX_BUSY,
        TX_DONE  => TX_DONE,
        RX       => RX,
        RX_BUSY  => RX_BUSY,
        RX_ERROR => RX_ERROR,
        RX_DATA  => RX_DATA
    );
--
PULSE_GEN : PROCESS(CLK)
  VARIABLE CNT_PULSE : INTEGER RANGE 0 TO 65535 := 0;
BEGIN
	IF CLK = '1' AND CLK'EVENT THEN
		IF CNT_PULSE < 4999 THEN
		    CNT_PULSE := CNT_PULSE + 1;
		ELSE 
		    CNT_PULSE := 0;
		END IF;
		IF CNT_PULSE < 100 THEN
			PULSE <= '1';
		ELSE
			PULSE <= '0';
		END IF;
	END IF;
END PROCESS;
--
RST_GEN : PROCESS(CLK)
  VARIABLE CNT_RST : INTEGER RANGE 0 TO 10000000 := 0;
BEGIN
	IF CLK = '1' AND CLK'EVENT THEN
		IF CNT_RST < 10000000 THEN
		    CNT_RST := CNT_RST + 1;
		ELSE 
		    CNT_RST := 0;
		END IF;
		IF CNT_RST < 20000 THEN
			RST_N <= '0';
		ELSE
			RST_N <= '1';
		END IF;
	END IF;
END PROCESS;
--
TRAN_GEN: PROCESS(CLK, RST_N)
BEGIN
    IF RST_N = '0' THEN
        TX_ENA <= '0';
        CNT_DATA <= X"0000";
    ELSIF rising_edge(CLK) THEN
        TX_ENA <= '0';
        IF CNT_DATA < X"0006" THEN
            TX_ENA <= PULSE;
            TX_DATA <= HELLO(CONV_INTEGER(CNT_DATA));
        END IF;
        IF TX_DONE = '1' THEN
            CNT_DATA <= CNT_DATA + X"0001";
            IF CNT_DATA = X"000A" THEN
                CNT_DATA <= X"0000";
            END IF;
        END IF;
    END IF;
END PROCESS;


END TRANSFER_ARCH;	
